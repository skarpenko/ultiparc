/*
 * Copyright (c) 2015-2016 The Ultiparc Project. All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
 * OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
 * LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */

/*
 * Register names
 */


/* General purpose registers */
localparam [4:0] R0  = 5'd0;
localparam [4:0] R1  = 5'd1;
localparam [4:0] R2  = 5'd2;
localparam [4:0] R3  = 5'd3;
localparam [4:0] R4  = 5'd4;
localparam [4:0] R5  = 5'd5;
localparam [4:0] R6  = 5'd6;
localparam [4:0] R7  = 5'd7;
localparam [4:0] R8  = 5'd8;
localparam [4:0] R9  = 5'd9;
localparam [4:0] R10 = 5'd10;
localparam [4:0] R11 = 5'd11;
localparam [4:0] R12 = 5'd12;
localparam [4:0] R13 = 5'd13;
localparam [4:0] R14 = 5'd14;
localparam [4:0] R15 = 5'd15;
localparam [4:0] R16 = 5'd16;
localparam [4:0] R17 = 5'd17;
localparam [4:0] R18 = 5'd18;
localparam [4:0] R19 = 5'd19;
localparam [4:0] R20 = 5'd20;
localparam [4:0] R21 = 5'd21;
localparam [4:0] R22 = 5'd22;
localparam [4:0] R23 = 5'd23;
localparam [4:0] R24 = 5'd24;
localparam [4:0] R25 = 5'd25;
localparam [4:0] R26 = 5'd26;
localparam [4:0] R27 = 5'd27;
localparam [4:0] R28 = 5'd28;
localparam [4:0] R29 = 5'd29;
localparam [4:0] R30 = 5'd30;
localparam [4:0] R31 = 5'd31;
