/*
 * Copyright (c) 2015-2016 The Ultiparc Project. All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
 * OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
 * LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */

/*
 * Fabric port FSM
 */

`include "common.vh"
`include "ocp_const.vh"


/*
 * Fabric port FSM
 */
module fabric_port #(
	parameter [10:0] PORT = 0	/* Port number */
)
(
	clk,
	nrst,
	/* OCP interface: instructions (master) */
	i_I_MAddr,
	i_I_MCmd,
	i_I_MData,
	i_I_MByteEn,
	o_I_SCmdAccept,
	o_I_SData,
	o_I_SResp,
	/* OCP interface: data (master) */
	i_D_MAddr,
	i_D_MCmd,
	i_D_MData,
	i_D_MByteEn,
	o_D_SCmdAccept,
	o_D_SData,
	o_D_SResp,
	/* OCP interface: Port (slave) */
	o_P_MAddr,
	o_P_MCmd,
	o_P_MData,
	o_P_MByteEn,
	i_P_SCmdAccept,
	i_P_SData,
	i_P_SResp
);
localparam PORT_BITS = 12;

input wire			clk;
input wire			nrst;
/* OCP interface: instructions */
input wire [`ADDR_WIDTH-1:0]	i_I_MAddr;
input wire [2:0]		i_I_MCmd;
input wire [`DATA_WIDTH-1:0]	i_I_MData;
input wire [`BEN_WIDTH-1:0]	i_I_MByteEn;
output wire			o_I_SCmdAccept;
output wire [`DATA_WIDTH-1:0]	o_I_SData;
output wire [1:0]		o_I_SResp;
/* OCP interface: data */
input wire [`ADDR_WIDTH-1:0]	i_D_MAddr;
input wire [2:0]		i_D_MCmd;
input wire [`DATA_WIDTH-1:0]	i_D_MData;
input wire [`BEN_WIDTH-1:0]	i_D_MByteEn;
output wire			o_D_SCmdAccept;
output wire [`DATA_WIDTH-1:0]	o_D_SData;
output wire [1:0]		o_D_SResp;
/* OCP interface: Port */
output wire [`ADDR_WIDTH-1:0]	o_P_MAddr;
output wire [2:0]		o_P_MCmd;
output wire [`DATA_WIDTH-1:0]	o_P_MData;
output wire [`BEN_WIDTH-1:0]	o_P_MByteEn;
input wire			i_P_SCmdAccept;
input wire [`DATA_WIDTH-1:0]	i_P_SData;
input wire [1:0]		i_P_SResp;


/* Bus interface FSM states */
localparam [4:0] IDLE   = 5'b00001;	/* Idle state */
localparam [4:0] RUN    = 5'b00010;	/* Start transaction */
localparam [4:0] DWAIT  = 5'b00100;	/* Wait for slave data */
localparam [4:0] CWAIT  = 5'b01000;	/* Conflict wait */
localparam [4:0] BWAIT  = 5'b10000;	/* Wait for bus ready */


/* Bus FSM state */
reg [6:0] i_bus_state;
reg [6:0] i_bus_next_state;
reg [6:0] d_bus_state;
reg [6:0] d_bus_next_state;


/* Command accept signals */
assign o_I_SCmdAccept = ((i_bus_state == IDLE || i_I_MCmd == `OCP_CMD_IDLE) ? 1'b1 : 1'b0);
assign o_D_SCmdAccept = ((d_bus_state == IDLE || i_D_MCmd == `OCP_CMD_IDLE) ? 1'b1 : 1'b0);


/* Return port number */
function [PORT_BITS-2:0] port_no;
	input [`ADDR_WIDTH-1:0] addr;
	port_no = (addr[`ADDR_WIDTH-1] ? addr[`ADDR_WIDTH-2:`ADDR_WIDTH-PORT_BITS] + 1 : 0);
endfunction


/* Decode address */
function [`ADDR_WIDTH-1:0] decode_addr;
	input [`ADDR_WIDTH-1:0] addr;
	decode_addr = (!addr[`ADDR_WIDTH-1] ? { 1'b0, addr[`ADDR_WIDTH-2:0] } :
		{ {(PORT_BITS){1'b0}}, addr[`ADDR_WIDTH-PORT_BITS-1:0] });
endfunction


/* Check for conflict */
function confl;
	input [`ADDR_WIDTH-1:0] i_addr;
	input [2:0] i_cmd;
	input [`ADDR_WIDTH-1:0] d_addr;
	input [2:0] d_cmd;
	confl = (port_no(i_addr) == port_no(d_addr) &&
		i_cmd != `OCP_CMD_IDLE && d_cmd != `OCP_CMD_IDLE);
endfunction


/* Latched instructions port inputs */
reg [`ADDR_WIDTH-1:0]		i_addr;
reg [2:0]			i_cmd;
reg [`DATA_WIDTH-1:0]		i_data;
reg [`BEN_WIDTH-1:0]		i_ben;

/* Latched data port inputs */
reg [`ADDR_WIDTH-1:0]		d_addr;
reg [2:0]			d_cmd;
reg [`DATA_WIDTH-1:0]		d_data;
reg [`BEN_WIDTH-1:0]		d_ben;

/* Internal instructions port connections */
reg [`ADDR_WIDTH-1:0]		I_MAddr;
reg [2:0]			I_MCmd;
reg [`DATA_WIDTH-1:0]		I_MData;
reg [`BEN_WIDTH-1:0]		I_MByteEn;
wire [`DATA_WIDTH-1:0]		I_SData;
wire [1:0]			I_SResp;
wire				I_SCmdAccept;

/* Internal data port connections */
reg [`ADDR_WIDTH-1:0]		D_MAddr;
reg [2:0]			D_MCmd;
reg [`DATA_WIDTH-1:0]		D_MData;
reg [`BEN_WIDTH-1:0]		D_MByteEn;
wire [`DATA_WIDTH-1:0]		D_SData;
wire [1:0]			D_SResp;
wire				D_SCmdAccept;


reg i_busy;	/* Instruction fetch on the fly */
reg d_busy;	/* Data fetch on the fly */

wire select;

assign select = (d_busy ? 1'b0 : 1'b1);	/* Select port */


/* Force outputs to zero if in idle state */
assign o_I_SData = I_SData & (i_bus_state == IDLE ? {(`DATA_WIDTH){1'b0}} :
	{(`DATA_WIDTH){1'b1}} );
assign o_I_SResp = I_SResp & (i_bus_state == IDLE ? 2'b00 : 2'b11 );
assign o_D_SData = D_SData & (d_bus_state == IDLE ? {(`DATA_WIDTH){1'b0}} :
	{(`DATA_WIDTH){1'b1}} );
assign o_D_SResp = D_SResp & (d_bus_state == IDLE ? 2'b00 : 2'b11 );


/* Latch inputs */
always @(posedge clk)
begin
	i_addr <= i_I_MAddr;
	i_cmd <= i_I_MCmd;
	i_data <= i_I_MData;
	i_ben <= i_I_MByteEn;
	d_addr <= i_D_MAddr;
	d_cmd <= i_D_MCmd;
	d_data <= i_D_MData;
	d_ben <= i_D_MByteEn;
end


/* Seq logic */
always @(posedge clk or negedge nrst)
begin
	i_bus_state <= nrst ? i_bus_next_state : IDLE;
	d_bus_state <= nrst ? d_bus_next_state : IDLE;
end


/* Next state logic for instructions port */
always @(*)
begin : instructions_port
	i_bus_next_state = IDLE;

	if(i_bus_state == IDLE && i_I_MCmd != `OCP_CMD_IDLE && port_no(i_I_MAddr) == PORT)
		i_bus_next_state = RUN;
	else if(i_bus_state == RUN && (confl(i_I_MAddr, i_I_MCmd, i_D_MAddr, i_D_MCmd) || d_busy || !i_busy))
		i_bus_next_state = CWAIT;
	else if(i_bus_state == RUN && I_SCmdAccept == 1'b0)
		i_bus_next_state = BWAIT;
	else if(i_bus_state == RUN)
		i_bus_next_state = DWAIT;
	else if(i_bus_state == CWAIT && !d_busy && i_busy && I_SCmdAccept == 1'b0)
		i_bus_next_state = BWAIT;
	else if(i_bus_state == CWAIT && !d_busy && i_busy)
		i_bus_next_state = DWAIT;
	else if(i_bus_state == CWAIT)
		i_bus_next_state = CWAIT;
	else if(i_bus_state == BWAIT && I_SCmdAccept == 1'b0)
		i_bus_next_state = BWAIT;
	else if(i_bus_state == BWAIT && i_P_SResp != `OCP_RESP_NULL)
		i_bus_next_state = IDLE;
	else if(i_bus_state == BWAIT)
		i_bus_next_state = DWAIT;
	else if(i_bus_state == DWAIT && i_P_SResp != `OCP_RESP_NULL)
		i_bus_next_state = IDLE;
	else if(i_bus_state == DWAIT)
		i_bus_next_state = DWAIT;
end


/* Next state logic for data port */
always @(*)
begin : data_port
	d_bus_next_state = IDLE;

	if(d_bus_state == IDLE && i_D_MCmd != `OCP_CMD_IDLE && port_no(i_D_MAddr) == PORT)
		d_bus_next_state = RUN;
	else if(d_bus_state == RUN && (i_busy || !d_busy))
		d_bus_next_state = CWAIT;
	else if(d_bus_state == RUN && D_SCmdAccept == 1'b0)
		d_bus_next_state = BWAIT;
	else if(d_bus_state == RUN)
		d_bus_next_state = DWAIT;
	else if(d_bus_state == CWAIT && !i_busy && d_busy && D_SCmdAccept == 1'b0)
		d_bus_next_state = BWAIT;
	else if(d_bus_state == CWAIT && !i_busy && d_busy)
		d_bus_next_state = DWAIT;
	else if(d_bus_state == CWAIT)
		d_bus_next_state = CWAIT;
	else if(d_bus_state == BWAIT && D_SCmdAccept == 1'b0)
		d_bus_next_state = BWAIT;
	else if(d_bus_state == BWAIT && i_P_SResp != `OCP_RESP_NULL)
		d_bus_next_state = IDLE;
	else if(d_bus_state == BWAIT)
		d_bus_next_state = DWAIT;
	else if(d_bus_state == DWAIT && i_P_SResp != `OCP_RESP_NULL)
		d_bus_next_state = IDLE;
	else if(d_bus_state == DWAIT)
		d_bus_next_state = DWAIT;
end


/* Output logic for instructions port */
always @(i_bus_state or d_busy)
begin
	if(i_bus_state == IDLE)
	begin
		I_MAddr <= {(`ADDR_WIDTH){1'b0}};
		I_MCmd <= 3'b0;
		I_MData <= {(`DATA_WIDTH){1'b0}};
		I_MByteEn <= {(`BEN_WIDTH){1'b0}};
		i_busy <= 1'b0;
	end
	else if(i_bus_state == RUN)
	begin
		I_MAddr <= decode_addr(i_addr);
		I_MCmd <= i_cmd;
		I_MData <= i_data;
		I_MByteEn <= i_ben;
		if(!confl(i_addr, i_cmd, d_addr, d_cmd) && !d_busy)
			i_busy <= 1'b1;
	end
	else if(i_bus_state == CWAIT)
	begin
		i_busy <= (!d_busy ? 1'b1 : 1'b0);
	end
	else if(i_bus_state == DWAIT)
	begin
		I_MAddr <= {(`ADDR_WIDTH){1'b0}};
		I_MCmd <= 3'b0;
		I_MData <= {(`DATA_WIDTH){1'b0}};
		I_MByteEn <= {(`BEN_WIDTH){1'b0}};
	end
end


/* Output logic for data port */
always @(d_bus_state or i_busy)
begin
	if(d_bus_state == IDLE)
	begin
		D_MAddr <= {(`ADDR_WIDTH){1'b0}};
		D_MCmd <= 3'b0;
		D_MData <= {(`DATA_WIDTH){1'b0}};
		D_MByteEn <= {(`BEN_WIDTH){1'b0}};
		d_busy <= 1'b0;
	end
	else if(d_bus_state == RUN)
	begin
		D_MAddr <= decode_addr(d_addr);
		D_MCmd <= d_cmd;
		D_MData <= d_data;
		D_MByteEn <= d_ben;
		if(!i_busy)
			d_busy <= 1'b1;
	end
	else if(d_bus_state == CWAIT)
	begin
		d_busy <= (!i_busy ? 1'b1 : 1'b0);
	end
	else if(d_bus_state == DWAIT)
	begin
		D_MAddr <= {(`ADDR_WIDTH){1'b0}};
		D_MCmd <= 3'b0;
		D_MData <= {(`DATA_WIDTH){1'b0}};
		D_MByteEn <= {(`BEN_WIDTH){1'b0}};
	end
end


/* Ports demultiplexer */
fabric_port_demux demux(
	.i_select(select),
	.i_I_MAddr(I_MAddr),
	.i_I_MCmd(I_MCmd),
	.i_I_MData(I_MData),
	.i_I_MByteEn(I_MByteEn),
	.o_I_SCmdAccept(I_SCmdAccept),
	.o_I_SData(I_SData),
	.o_I_SResp(I_SResp),
	.i_D_MAddr(D_MAddr),
	.i_D_MCmd(D_MCmd),
	.i_D_MData(D_MData),
	.i_D_MByteEn(D_MByteEn),
	.o_D_SCmdAccept(D_SCmdAccept),
	.o_D_SData(D_SData),
	.o_D_SResp(D_SResp),
	.o_P_MAddr(o_P_MAddr),
	.o_P_MCmd(o_P_MCmd),
	.o_P_MData(o_P_MData),
	.o_P_MByteEn(o_P_MByteEn),
	.i_P_SCmdAccept(i_P_SCmdAccept),
	.i_P_SData(i_P_SData),
	.i_P_SResp(i_P_SResp)
);


endmodule /* fabric_port */
