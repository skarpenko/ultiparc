module cpu_top();
endmodule /* cpu_top */
